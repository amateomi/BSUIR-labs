module dist_arithmetic(
    input clk,
    input reset,
    input [7:0] x_msb,
    input [7:0] x_lsb,
    output [16:0] y,
    output valid
);

integer counter = 0;
always @(posedge clk or negedge reset)
begin
    if (reset)
        counter <= 0;
    else
        counter <= counter + 1;
end

reg signed [16:0] acc = 0;
assign valid = counter == 8;
assign y = valid ? acc : 0;

reg signed [16:0] ROM[127:0];
initial begin
    ROM[0] =   17'b11110100000000000;
    ROM[1] =   17'b11100100000000000;
    ROM[2] =   17'b11111100000000000;
    ROM[3] =   17'b11101100000000000;
    ROM[4] =   17'b11010100000000000;
    ROM[5] =   17'b11000100000000000;
    ROM[6] =   17'b11011100000000000;
    ROM[7] =   17'b11001100000000000;
    ROM[8] =   17'b00011100000000000;
    ROM[9] =   17'b00001100000000000;
    ROM[10] =  17'b00100100000000000;
    ROM[11] =  17'b00010100000000000;
    ROM[12] =  17'b11111100000000000;
    ROM[13] =  17'b11101100000000000;
    ROM[14] =  17'b00000100000000000;
    ROM[15] =  17'b11110100000000000;
    ROM[16] =  17'b11100100000000000;
    ROM[17] =  17'b11010100000000000;
    ROM[18] =  17'b11101100000000000;
    ROM[19] =  17'b11011100000000000;
    ROM[20] =  17'b11000100000000000;
    ROM[21] =  17'b10110100000000000;
    ROM[22] =  17'b11001100000000000;
    ROM[23] =  17'b10111100000000000;
    ROM[24] =  17'b00001100000000000;
    ROM[25] =  17'b11111100000000000;
    ROM[26] =  17'b00010100000000000;
    ROM[27] =  17'b00000100000000000;
    ROM[28] =  17'b11101100000000000;
    ROM[29] =  17'b11011100000000000;
    ROM[30] =  17'b11110100000000000;
    ROM[31] =  17'b11100100000000000;
    ROM[32] =  17'b11111100000000000;
    ROM[33] =  17'b11101100000000000;
    ROM[34] =  17'b00000100000000000;
    ROM[35] =  17'b11110100000000000;
    ROM[36] =  17'b11011100000000000;
    ROM[37] =  17'b11001100000000000;
    ROM[38] =  17'b11100100000000000;
    ROM[39] =  17'b11010100000000000;
    ROM[40] =  17'b00100100000000000;
    ROM[41] =  17'b00010100000000000;
    ROM[42] =  17'b00101100000000000;
    ROM[43] =  17'b00011100000000000;
    ROM[44] =  17'b00000100000000000;
    ROM[45] =  17'b11110100000000000;
    ROM[46] =  17'b00001100000000000;
    ROM[47] =  17'b11111100000000000;
    ROM[48] =  17'b11101100000000000;
    ROM[49] =  17'b11011100000000000;
    ROM[50] =  17'b11110100000000000;
    ROM[51] =  17'b11100100000000000;
    ROM[52] =  17'b11001100000000000;
    ROM[53] =  17'b10111100000000000;
    ROM[54] =  17'b11010100000000000;
    ROM[55] =  17'b11000100000000000;
    ROM[56] =  17'b00010100000000000;
    ROM[57] =  17'b00000100000000000;
    ROM[58] =  17'b00011100000000000;
    ROM[59] =  17'b00001100000000000;
    ROM[60] =  17'b11110100000000000;
    ROM[61] =  17'b11100100000000000;
    ROM[62] =  17'b11111100000000000;
    ROM[63] =  17'b11101100000000000;
    ROM[64] =  17'b00000100000000000;
    ROM[65] =  17'b11110100000000000;
    ROM[66] =  17'b00001100000000000;
    ROM[67] =  17'b11111100000000000;
    ROM[68] =  17'b11100100000000000;
    ROM[69] =  17'b11010100000000000;
    ROM[70] =  17'b11101100000000000;
    ROM[71] =  17'b11011100000000000;
    ROM[72] =  17'b00101100000000000;
    ROM[73] =  17'b00011100000000000;
    ROM[74] =  17'b00110100000000000;
    ROM[75] =  17'b00100100000000000;
    ROM[76] =  17'b00001100000000000;
    ROM[77] =  17'b11111100000000000;
    ROM[78] =  17'b00010100000000000;
    ROM[79] =  17'b00000100000000000;
    ROM[80] =  17'b11110100000000000;
    ROM[81] =  17'b11100100000000000;
    ROM[82] =  17'b11111100000000000;
    ROM[83] =  17'b11101100000000000;
    ROM[84] =  17'b11010100000000000;
    ROM[85] =  17'b11000100000000000;
    ROM[86] =  17'b11011100000000000;
    ROM[87] =  17'b11001100000000000;
    ROM[88] =  17'b00011100000000000;
    ROM[89] =  17'b00001100000000000;
    ROM[90] =  17'b00100100000000000;
    ROM[91] =  17'b00010100000000000;
    ROM[92] =  17'b11111100000000000;
    ROM[93] =  17'b11101100000000000;
    ROM[94] =  17'b00000100000000000;
    ROM[95] =  17'b11110100000000000;
    ROM[96] =  17'b00001100000000000;
    ROM[97] =  17'b11111100000000000;
    ROM[98] =  17'b00010100000000000;
    ROM[99] =  17'b00000100000000000;
    ROM[100] = 17'b11101100000000000;
    ROM[101] = 17'b11011100000000000;
    ROM[102] = 17'b11110100000000000;
    ROM[103] = 17'b11100100000000000;
    ROM[104] = 17'b00110100000000000;
    ROM[105] = 17'b00100100000000000;
    ROM[106] = 17'b00111100000000000;
    ROM[107] = 17'b00101100000000000;
    ROM[108] = 17'b00010100000000000;
    ROM[109] = 17'b00000100000000000;
    ROM[110] = 17'b00011100000000000;
    ROM[111] = 17'b00001100000000000;
    ROM[112] = 17'b11111100000000000;
    ROM[113] = 17'b11101100000000000;
    ROM[114] = 17'b00000100000000000;
    ROM[115] = 17'b11110100000000000;
    ROM[116] = 17'b11011100000000000;
    ROM[117] = 17'b11001100000000000;
    ROM[118] = 17'b11100100000000000;
    ROM[119] = 17'b11010100000000000;
    ROM[120] = 17'b00100100000000000;
    ROM[121] = 17'b00010100000000000;
    ROM[122] = 17'b00101100000000000;
    ROM[123] = 17'b00011100000000000;
    ROM[124] = 17'b00000100000000000;
    ROM[125] = 17'b11110100000000000;
    ROM[126] = 17'b00001100000000000;
    ROM[127] = 17'b11111100000000000;
end

function [6:0] xored(input [7:0] x);
    begin
        xored = {x[7] ^ x[6],
                 x[7] ^ x[5],
                 x[7] ^ x[4],
                 x[7] ^ x[3],
                 x[7] ^ x[2],
                 x[7] ^ x[1],
                 x[7] ^ x[0]};
    end
endfunction

// Macro is used because the identical function does not work for some reason
`define fetch_from_ROM(x, ts) ((ts ^ x[7]) ? -ROM[xored(x)] : ROM[xored(x)])

always @(posedge clk or negedge reset)
begin
    if (reset)
        acc <= 0;
    else if (counter == 0)
        acc <= ((ROM[0] + `fetch_from_ROM(x_lsb, 0)) >>> 1) + `fetch_from_ROM(x_msb, 0);
    else if (counter == 7)
        acc <= (((acc >>> 1) + `fetch_from_ROM(x_lsb, 0)) >>> 1) + `fetch_from_ROM(x_msb, 1);
    else
        acc <= (((acc >>> 1) + `fetch_from_ROM(x_lsb, 0)) >>> 1) + `fetch_from_ROM(x_msb, 0);
end
endmodule
